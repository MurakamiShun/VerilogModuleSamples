`define FP_ROUND_TONEAREST  2'b00
`define FP_ROUND_TOWARDZERO 2'b01
`define FP_ROUND_DOWNWARD   2'b10
`define FP_ROUND_UPWARD     2'b11

// bit positions
`define FP_INVALID    4
`define FP_DIVBYZERO  3
`define FP_OVERFLOW   2
`define FP_UNDERFLOW  1
`define FP_INEXACT    0